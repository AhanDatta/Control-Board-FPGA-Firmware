module AD9228_core_testbench #(
    parameter DATA_WIDTH = 12
) ();

    

endmodule