//Take in cmnd from IPIF (AXI) interface
/*
Create IPIF struct with all values to be written
*/
//Update state machine
/*
detect new IPIF cmnd, by setting one of the bits as a self-reseting flag
Do cmnd
*/
//Send out command