//create writing state machine to send instructions
