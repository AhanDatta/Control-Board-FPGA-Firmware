module AD9228_core_emulator (
    input logic clk,
    input logic csb,

    output logic fco,
    output logic dco,
    output logic dout
);

    

endmodule